`ifndef __TABLE_LOGGER_PKG_SV__
`define __TABLE_LOGGER_PKG_SV__

package table_logger_pkg;

  import uvm_pkg::*;
  `include "uvm_macros.svh"

  `include "txt_tbl.sv"
  `include "enum_width_finder.svh"
  `include "table_logger_cfg.svh"
  `include "table_logger.svh"

endpackage

`endif
