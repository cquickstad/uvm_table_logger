typedef enum bit [1:0] {
    FIRST_ENUM_VALUE,
    SECOND_ENUM_VALUE,
    THIRD_ENUM_VALUE,
    LAST_ENUM_VALUE
} my_enum_t;
