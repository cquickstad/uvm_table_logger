// -------------------------------------------------------------
//    Copyright 2020 Chad Quickstad
//    All Rights Reserved Worldwide
//
//    Licensed under the Apache License, Version 2.0 (the
//    "License"); you may not use this file except in
//    compliance with the License.  You may obtain a copy of
//    the License at
//
//        http://www.apache.org/licenses/LICENSE-2.0
//
//    Unless required by applicable law or agreed to in
//    writing, software distributed under the License is
//    distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
//    CONDITIONS OF ANY KIND, either express or implied.  See
//    the License for the specific language governing
//    permissions and limitations under the License.
// -------------------------------------------------------------

// Look for the latest version of this code at:
//  https://github.com/cquickstad/uvm_table_logger.git

`ifndef __MY_PKG_SV__
`define __MY_PKG_SV__

package my_pkg;

  import uvm_pkg::*;
  `include "uvm_macros.svh"

  `include "my_types.svh"
  `include "my_item.svh"
  `include "my_sequencer.svh"
  `include "my_driver.svh"
  `include "my_monitor.svh"
  `include "my_agent.svh"
  `include "my_table_item.svh"
  `include "my_env.svh"
  `include "my_sequence_base.svh"
  `include "my_sequence_lib.svh"
  `include "my_vseq_base.svh"
  `include "my_vseq_lib.svh"
  `include "my_test_base.svh"
  `include "my_test_lib.svh"

endpackage

`endif
